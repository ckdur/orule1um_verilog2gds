VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.25 ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

# High density, single height
SITE obscore
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 2.0 BY 40.0 ;
END obscore

#--------EOF---------

MACRO AN2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1 0 0 ; 
  SIZE 28.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 20.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 0.000 39.000 28.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 28.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 0.000 -1.000 28.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 28.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 6.500 14.250 21.500 ;
        RECT 12.750 20.000 14.750 22.000 ;
  END
END AN2D1
MACRO AN2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1_1 0 0 ; 
  SIZE 22.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a2 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 20.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 0.000 39.000 22.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 22.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.000 -1.000 22.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 22.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 1.250 6.500 11.250 7.500 ;
        RECT 10.250 2.500 11.250 7.500 ;
        RECT 9.750 2.000 11.750 4.000 ;
        RECT 7.250 6.500 8.250 30.500 ;
  END
END AN2D1_1
MACRO AN2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1_2 0 0 ; 
  SIZE 28.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 20.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 0.000 39.000 28.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 28.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 0.000 -1.000 28.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 28.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 6.500 14.250 21.500 ;
        RECT 12.750 20.000 14.750 22.000 ;
  END
END AN2D1_2
MACRO AN2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AN2D1_3 0 0 ; 
  SIZE 28.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a2 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 20.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 0.000 39.000 28.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 28.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.000 -1.000 28.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 28.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 1.250 6.500 2.250 25.500 ;
        RECT 1.250 24.500 14.250 25.500 ;
        RECT 13.250 24.500 14.250 30.500 ;
  END
END AN2D1_3
#--------EOF---------

MACRO AO21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1 0 0 ; 
  SIZE 34.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END b 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 6.500 26.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 29.500 32.250 39.500 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 29.500 20.250 39.500 ;
        RECT 0.000 39.000 34.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 34.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 31.250 0.500 32.250 7.500 ;
        RECT 0.000 -1.000 34.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 34.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 1.250 2.500 2.250 7.500 ;
        RECT 0.750 2.000 2.750 4.000 ;
        RECT 19.250 2.500 20.250 7.500 ;
        RECT 19.250 2.500 29.250 3.500 ;
        RECT 27.750 2.000 29.750 4.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 1.250 29.500 14.250 30.500 ;
  END
END AO21D1
MACRO AO21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1_1 0 0 ; 
  SIZE 34.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 22.250 14.500 23.250 18.500 ;
    END 
  END b 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 6.500 32.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 0.000 39.000 34.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 34.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 0.000 -1.000 34.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 34.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 2.500 14.250 7.500 ;
        RECT 12.750 2.000 14.750 4.000 ;
        RECT 15.750 29.000 17.750 31.000 ;
        RECT 13.250 29.500 17.250 30.500 ;
        RECT 16.250 6.500 20.250 7.500 ;
        RECT 15.750 6.000 17.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 7.250 24.500 8.250 30.500 ;
        RECT 7.250 24.500 20.250 25.500 ;
        RECT 19.250 24.500 20.250 30.500 ;
  END
END AO21D1_1
MACRO AO21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1_2 0 0 ; 
  SIZE 34.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END b 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 6.500 26.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 29.500 32.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 0.000 39.000 34.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 34.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 31.250 0.500 32.250 7.500 ;
        RECT 0.000 -1.000 34.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 34.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 7.250 6.500 8.250 25.500 ;
        RECT 7.250 24.500 14.250 25.500 ;
        RECT 13.250 24.500 14.250 30.500 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 7.250 29.500 8.250 33.500 ;
        RECT 7.250 32.500 20.250 33.500 ;
        RECT 19.250 29.500 20.250 33.500 ;
  END
END AO21D1_2
MACRO AO21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21D1_3 0 0 ; 
  SIZE 34.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END b 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 6.500 26.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 29.500 32.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 0.000 39.000 34.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 34.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 31.250 0.500 32.250 7.500 ;
        RECT 0.000 -1.000 34.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 34.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 19.250 2.500 20.250 7.500 ;
        RECT 19.250 2.500 29.250 3.500 ;
        RECT 27.750 2.000 29.750 4.000 ;
        RECT 1.250 2.500 2.250 7.500 ;
        RECT 0.750 2.000 2.750 4.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 20.250 30.500 ;
  END
END AO21D1_3
#--------EOF---------

MACRO AOI21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1 0 0 ; 
  SIZE 22.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END b 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 13.250 6.500 14.250 25.500 ;
        RECT 7.250 24.500 14.250 25.500 ;
        RECT 7.250 24.500 8.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 29.500 20.250 39.500 ;
        RECT 0.000 39.000 22.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 22.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 0.000 -1.000 22.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 22.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 1.250 29.500 2.250 33.500 ;
        RECT 1.250 32.500 14.250 33.500 ;
        RECT 13.250 29.500 14.250 33.500 ;
  END
END AOI21D1
MACRO AOI21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1_1 0 0 ; 
  SIZE 22.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END b 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 7.250 6.500 8.250 25.500 ;
        RECT 7.250 24.500 14.250 25.500 ;
        RECT 13.250 24.500 14.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 0.000 39.000 22.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 22.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 0.000 -1.000 22.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 22.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 19.250 29.500 20.250 33.500 ;
        RECT 7.250 32.500 20.250 33.500 ;
        RECT 7.250 29.500 8.250 33.500 ;
  END
END AOI21D1_1
MACRO AOI21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1_2 0 0 ; 
  SIZE 28.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 14.000 2.750 16.000 ;
        RECT 1.250 14.500 2.250 18.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 22.250 14.500 23.250 18.500 ;
    END 
  END b 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 4.250 6.500 14.250 7.500 ;
        RECT 4.250 6.500 5.250 30.500 ;
        RECT 1.250 29.500 5.250 30.500 ;
        RECT 13.250 6.500 20.250 7.500 ;
        RECT 4.250 29.500 5.250 33.500 ;
        RECT 4.250 32.500 14.250 33.500 ;
        RECT 13.250 29.500 14.250 33.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 0.000 39.000 28.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 28.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 0.000 -1.000 28.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 28.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 7.250 24.500 8.250 30.500 ;
        RECT 7.250 24.500 20.250 25.500 ;
        RECT 19.250 24.500 20.250 30.500 ;
  END
END AOI21D1_2
MACRO AOI21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21D1_3 0 0 ; 
  SIZE 28.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 22.250 14.500 23.250 18.500 ;
    END 
  END b 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 6.500 2.250 30.500 ;
        RECT 19.250 6.500 20.250 25.500 ;
        RECT 13.250 24.500 20.250 25.500 ;
        RECT 13.250 24.500 14.250 30.500 ;
        RECT 1.250 24.500 14.250 25.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 0.000 39.000 28.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 28.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 0.000 -1.000 28.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 28.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 7.250 29.500 8.250 33.500 ;
        RECT 7.250 32.500 20.250 33.500 ;
        RECT 19.250 29.500 20.250 33.500 ;
  END
END AOI21D1_3
#--------EOF---------

MACRO BUFFD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFFD1 0 0 ; 
  SIZE 16.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN i 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 17.000 11.750 19.000 ;
        RECT 10.250 17.500 11.250 25.500 ;
        RECT 9.750 24.000 11.750 26.000 ;
    END 
  END i 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 6.500 2.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 0.000 39.000 16.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 16.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 0.000 -1.000 16.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 16.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 12.750 24.000 14.750 26.000 ;
        RECT 13.250 24.500 14.250 30.500 ;
        RECT 13.250 6.500 14.250 21.500 ;
        RECT 12.750 20.000 14.750 22.000 ;
  END
END BUFFD1
MACRO BUFFD1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFFD1_1 0 0 ; 
  SIZE 16.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN i 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END i 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 6.500 14.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 0.000 39.000 16.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 16.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 0.000 -1.000 16.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 16.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 6.500 2.250 30.500 ;
  END
END BUFFD1_1
#--------EOF---------

MACRO DFCNQD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFCNQD1 0 0 ; 
  SIZE 106.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN cdn 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 45.750 2.000 47.750 4.000 ;
        RECT 43.250 2.500 47.250 3.500 ;
    END 
  END cdn 
  PIN cp 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END cp 
  PIN d 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 14.000 26.750 16.000 ;
        RECT 25.250 14.500 26.250 18.500 ;
    END 
  END d 
  PIN q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 102.750 6.000 104.750 8.000 ;
        RECT 96.750 29.000 98.750 31.000 ;
        RECT 103.250 6.500 104.250 25.500 ;
        RECT 97.250 24.500 104.250 25.500 ;
        RECT 97.250 24.500 98.250 30.500 ;
    END 
  END q 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 29.500 20.250 39.500 ;
        RECT 42.750 32.000 44.750 34.000 ;
        RECT 43.250 32.500 44.250 39.500 ;
        RECT 54.750 32.000 56.750 34.000 ;
        RECT 55.250 32.500 56.250 39.500 ;
        RECT 78.750 32.000 80.750 34.000 ;
        RECT 79.250 32.500 80.250 39.500 ;
        RECT 90.750 29.000 92.750 31.000 ;
        RECT 91.250 29.500 92.250 39.500 ;
        RECT 0.000 39.000 106.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 106.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 48.750 6.000 50.750 8.000 ;
        RECT 49.250 0.500 50.250 7.500 ;
        RECT 78.750 6.000 80.750 8.000 ;
        RECT 79.250 0.500 80.250 7.500 ;
        RECT 96.750 6.000 98.750 8.000 ;
        RECT 97.250 0.500 98.250 7.500 ;
        RECT 0.000 -1.000 106.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 106.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 6.500 5.250 7.500 ;
        RECT 4.250 2.500 5.250 7.500 ;
        RECT 3.750 2.000 5.750 4.000 ;
        RECT 1.250 6.500 2.250 30.500 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 6.500 17.250 7.500 ;
        RECT 16.250 6.500 17.250 11.500 ;
        RECT 16.250 10.500 29.250 11.500 ;
        RECT 28.250 2.500 29.250 11.500 ;
        RECT 28.250 2.500 35.250 3.500 ;
        RECT 33.750 2.000 35.750 4.000 ;
        RECT 28.250 10.500 29.250 37.500 ;
        RECT 28.250 36.500 41.250 37.500 ;
        RECT 39.750 36.000 41.750 38.000 ;
        RECT 63.750 36.000 65.750 38.000 ;
        RECT 64.250 14.500 65.250 37.500 ;
        RECT 58.250 14.500 65.250 15.500 ;
        RECT 57.750 14.000 59.750 16.000 ;
        RECT 13.250 6.500 14.250 30.500 ;
        RECT 22.250 20.500 29.250 21.500 ;
        RECT 21.750 20.000 23.750 22.000 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 6.500 47.250 7.500 ;
        RECT 46.250 6.500 47.250 15.500 ;
        RECT 46.250 14.500 53.250 15.500 ;
        RECT 51.750 14.000 53.750 16.000 ;
        RECT 31.250 6.500 32.250 30.500 ;
        RECT 36.750 32.000 38.750 34.000 ;
        RECT 48.750 32.000 50.750 34.000 ;
        RECT 37.250 32.500 41.250 33.500 ;
        RECT 40.250 29.500 41.250 33.500 ;
        RECT 40.250 29.500 50.250 30.500 ;
        RECT 49.250 29.500 50.250 33.500 ;
        RECT 54.750 6.000 56.750 8.000 ;
        RECT 60.750 29.000 62.750 31.000 ;
        RECT 39.750 14.000 41.750 16.000 ;
        RECT 40.250 14.500 44.250 15.500 ;
        RECT 43.250 14.500 44.250 18.500 ;
        RECT 43.250 17.500 56.250 18.500 ;
        RECT 55.250 6.500 56.250 18.500 ;
        RECT 55.250 17.500 56.250 25.500 ;
        RECT 55.250 24.500 62.250 25.500 ;
        RECT 61.250 24.500 62.250 30.500 ;
        RECT 60.750 6.000 62.750 8.000 ;
        RECT 66.750 29.000 68.750 31.000 ;
        RECT 61.250 6.500 77.250 7.500 ;
        RECT 76.250 6.500 77.250 11.500 ;
        RECT 76.250 10.500 89.250 11.500 ;
        RECT 88.250 2.500 89.250 11.500 ;
        RECT 87.750 2.000 89.750 4.000 ;
        RECT 67.250 6.500 68.250 30.500 ;
        RECT 66.750 6.000 68.750 8.000 ;
        RECT 72.750 6.000 74.750 8.000 ;
        RECT 67.250 2.500 68.250 7.500 ;
        RECT 67.250 2.500 74.250 3.500 ;
        RECT 73.250 2.500 74.250 7.500 ;
        RECT 90.750 6.000 92.750 8.000 ;
        RECT 84.750 29.000 86.750 31.000 ;
        RECT 78.750 14.000 80.750 16.000 ;
        RECT 79.250 14.500 92.250 15.500 ;
        RECT 91.250 6.500 92.250 15.500 ;
        RECT 91.250 14.500 101.250 15.500 ;
        RECT 99.750 14.000 101.750 16.000 ;
        RECT 85.250 14.500 86.250 30.500 ;
        RECT 94.250 14.500 95.250 21.500 ;
        RECT 93.750 20.000 95.750 22.000 ;
  END
END DFCNQD1
#--------EOF---------

MACRO DFQD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1 0 0 ; 
  SIZE 94.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN cp 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END cp 
  PIN d 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END d 
  PIN q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 84.750 6.000 86.750 8.000 ;
        RECT 84.750 29.000 86.750 31.000 ;
        RECT 85.250 6.500 86.250 30.500 ;
    END 
  END q 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 32.000 32.750 34.000 ;
        RECT 31.250 32.500 32.250 39.500 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 90.750 29.000 92.750 31.000 ;
        RECT 91.250 29.500 92.250 39.500 ;
        RECT 54.750 29.000 56.750 31.000 ;
        RECT 55.250 29.500 56.250 39.500 ;
        RECT 66.750 32.000 68.750 34.000 ;
        RECT 67.250 32.500 68.250 39.500 ;
        RECT 0.000 39.000 94.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 94.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 31.250 0.500 32.250 7.500 ;
        RECT 66.750 6.000 68.750 8.000 ;
        RECT 67.250 0.500 68.250 7.500 ;
        RECT 90.750 6.000 92.750 8.000 ;
        RECT 91.250 0.500 92.250 7.500 ;
        RECT 54.750 6.000 56.750 8.000 ;
        RECT 55.250 0.500 56.250 7.500 ;
        RECT 0.000 -1.000 94.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 94.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 9.750 20.000 11.750 22.000 ;
        RECT 4.250 20.500 11.250 21.500 ;
        RECT 4.250 20.500 5.250 30.500 ;
        RECT 1.250 29.500 5.250 30.500 ;
        RECT 48.750 2.000 50.750 4.000 ;
        RECT 34.250 2.500 50.250 3.500 ;
        RECT 33.750 2.000 35.750 4.000 ;
        RECT 0.750 2.000 2.750 4.000 ;
        RECT 1.250 2.500 2.250 7.500 ;
        RECT 10.250 20.500 11.250 37.500 ;
        RECT 10.250 36.500 23.250 37.500 ;
        RECT 21.750 36.000 23.750 38.000 ;
        RECT 78.750 6.000 80.750 8.000 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 78.750 32.000 80.750 34.000 ;
        RECT 79.250 6.500 80.250 21.500 ;
        RECT 58.250 20.500 80.250 21.500 ;
        RECT 57.750 20.000 59.750 22.000 ;
        RECT 79.250 20.500 80.250 33.500 ;
        RECT 43.250 6.500 44.250 30.500 ;
        RECT 57.750 14.000 59.750 16.000 ;
        RECT 58.250 14.500 59.250 18.500 ;
        RECT 58.250 17.500 80.250 18.500 ;
        RECT 79.250 17.500 80.250 21.500 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 23.250 7.500 ;
        RECT 22.250 6.500 23.250 30.500 ;
        RECT 19.250 29.500 23.250 30.500 ;
        RECT 21.750 20.000 23.750 22.000 ;
        RECT 54.750 14.000 56.750 16.000 ;
        RECT 55.250 14.500 56.250 21.500 ;
        RECT 54.750 20.000 56.750 22.000 ;
        RECT 36.750 6.000 38.750 8.000 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 36.750 17.000 38.750 19.000 ;
        RECT 37.250 17.500 38.250 30.500 ;
        RECT 37.250 29.500 38.250 37.500 ;
        RECT 37.250 36.500 53.250 37.500 ;
        RECT 51.750 36.000 53.750 38.000 ;
        RECT 39.750 6.000 41.750 8.000 ;
        RECT 37.250 6.500 41.250 7.500 ;
        RECT 37.250 6.500 38.250 30.500 ;
        RECT 48.750 6.000 50.750 8.000 ;
        RECT 48.750 29.000 50.750 31.000 ;
        RECT 27.750 14.000 29.750 16.000 ;
        RECT 28.250 14.500 29.250 25.500 ;
        RECT 27.750 24.000 29.750 26.000 ;
        RECT 49.250 6.500 50.250 30.500 ;
        RECT 48.750 14.000 50.750 16.000 ;
        RECT 60.750 6.000 62.750 8.000 ;
        RECT 69.750 10.000 71.750 12.000 ;
        RECT 61.250 10.500 71.250 11.500 ;
        RECT 61.250 6.500 62.250 11.500 ;
  END
END DFQD1
MACRO DFQD1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1_1 0 0 ; 
  SIZE 88.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN cp 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 17.000 5.750 19.000 ;
        RECT 4.250 17.500 5.250 21.500 ;
    END 
  END cp 
  PIN d 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END d 
  PIN q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 78.750 6.000 80.750 8.000 ;
        RECT 78.750 29.000 80.750 31.000 ;
        RECT 79.250 6.500 80.250 30.500 ;
    END 
  END q 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 32.000 32.750 34.000 ;
        RECT 31.250 32.500 32.250 39.500 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 84.750 29.000 86.750 31.000 ;
        RECT 85.250 29.500 86.250 39.500 ;
        RECT 66.750 32.000 68.750 34.000 ;
        RECT 67.250 32.500 68.250 39.500 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 43.250 29.500 44.250 39.500 ;
        RECT 0.000 39.000 88.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 88.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 31.250 0.500 32.250 7.500 ;
        RECT 66.750 6.000 68.750 8.000 ;
        RECT 67.250 0.500 68.250 7.500 ;
        RECT 84.750 6.000 86.750 8.000 ;
        RECT 85.250 0.500 86.250 7.500 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 43.250 0.500 44.250 7.500 ;
        RECT 0.000 -1.000 88.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 88.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 1.250 14.500 11.250 15.500 ;
        RECT 1.250 14.500 2.250 30.500 ;
        RECT 1.250 29.500 2.250 37.500 ;
        RECT 0.750 36.000 2.750 38.000 ;
        RECT 1.250 6.500 2.250 15.500 ;
        RECT 54.750 6.000 56.750 8.000 ;
        RECT 54.750 29.000 56.750 31.000 ;
        RECT 55.250 2.500 56.250 7.500 ;
        RECT 54.750 2.000 56.750 4.000 ;
        RECT 55.250 6.500 62.250 7.500 ;
        RECT 61.250 6.500 62.250 18.500 ;
        RECT 61.250 17.500 71.250 18.500 ;
        RECT 69.750 17.000 71.750 19.000 ;
        RECT 61.250 17.500 62.250 25.500 ;
        RECT 55.250 24.500 62.250 25.500 ;
        RECT 55.250 24.500 56.250 30.500 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 18.750 32.000 20.750 34.000 ;
        RECT 19.250 6.500 20.250 30.500 ;
        RECT 19.250 32.500 26.250 33.500 ;
        RECT 25.250 32.500 26.250 37.500 ;
        RECT 24.750 36.000 26.750 38.000 ;
        RECT 36.750 6.000 38.750 8.000 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 21.750 24.000 23.750 26.000 ;
        RECT 22.250 24.500 23.250 30.500 ;
        RECT 22.250 29.500 38.250 30.500 ;
        RECT 21.750 17.000 23.750 19.000 ;
        RECT 22.250 17.500 59.250 18.500 ;
        RECT 57.750 17.000 59.750 19.000 ;
        RECT 36.750 2.000 38.750 4.000 ;
        RECT 37.250 2.500 38.250 7.500 ;
        RECT 51.750 17.000 53.750 19.000 ;
        RECT 48.750 6.000 50.750 8.000 ;
        RECT 48.750 29.000 50.750 31.000 ;
        RECT 27.750 10.000 29.750 12.000 ;
        RECT 28.250 10.500 50.250 11.500 ;
        RECT 49.250 6.500 50.250 11.500 ;
        RECT 49.250 10.500 50.250 15.500 ;
        RECT 48.750 14.000 50.750 16.000 ;
        RECT 48.750 20.000 50.750 22.000 ;
        RECT 49.250 20.500 50.250 30.500 ;
        RECT 28.250 24.500 50.250 25.500 ;
        RECT 27.750 24.000 29.750 26.000 ;
        RECT 72.750 6.000 74.750 8.000 ;
        RECT 63.750 10.000 65.750 12.000 ;
        RECT 64.250 10.500 71.250 11.500 ;
        RECT 70.250 2.500 71.250 11.500 ;
        RECT 70.250 2.500 83.250 3.500 ;
        RECT 81.750 2.000 83.750 4.000 ;
        RECT 70.250 6.500 74.250 7.500 ;
  END
END DFQD1_1
MACRO DFQD1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1_2 0 0 ; 
  SIZE 88.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN cp 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 10.500 5.250 15.500 ;
    END 
  END cp 
  PIN d 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 27.750 17.000 29.750 19.000 ;
        RECT 28.250 17.500 29.250 25.500 ;
        RECT 27.750 24.000 29.750 26.000 ;
    END 
  END d 
  PIN q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 78.750 6.000 80.750 8.000 ;
        RECT 78.750 29.000 80.750 31.000 ;
        RECT 76.250 6.500 80.250 7.500 ;
        RECT 75.750 6.000 77.750 8.000 ;
        RECT 75.750 29.000 77.750 31.000 ;
        RECT 76.250 29.500 80.250 30.500 ;
    END 
  END q 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 84.750 29.000 86.750 31.000 ;
        RECT 85.250 29.500 86.250 39.500 ;
        RECT 66.750 32.000 68.750 34.000 ;
        RECT 67.250 32.500 68.250 39.500 ;
        RECT 42.750 32.000 44.750 34.000 ;
        RECT 43.250 32.500 44.250 39.500 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 29.500 20.250 39.500 ;
        RECT 0.000 39.000 88.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 88.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 43.250 0.500 44.250 7.500 ;
        RECT 66.750 6.000 68.750 8.000 ;
        RECT 67.250 0.500 68.250 7.500 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 84.750 6.000 86.750 8.000 ;
        RECT 85.250 0.500 86.250 7.500 ;
        RECT 0.000 -1.000 88.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 88.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 57.750 10.000 59.750 12.000 ;
        RECT 58.250 10.500 59.250 18.500 ;
        RECT 52.250 17.500 59.250 18.500 ;
        RECT 51.750 17.000 53.750 19.000 ;
        RECT 3.750 17.000 5.750 19.000 ;
        RECT 4.250 17.500 5.250 30.500 ;
        RECT 1.250 29.500 5.250 30.500 ;
        RECT 1.250 6.500 2.250 18.500 ;
        RECT 1.250 17.500 8.250 18.500 ;
        RECT 6.750 17.000 8.750 19.000 ;
        RECT 1.250 17.500 5.250 18.500 ;
        RECT 54.750 6.000 56.750 8.000 ;
        RECT 54.750 32.000 56.750 34.000 ;
        RECT 55.250 2.500 56.250 7.500 ;
        RECT 54.750 2.000 56.750 4.000 ;
        RECT 54.750 36.000 56.750 38.000 ;
        RECT 55.250 32.500 56.250 37.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 6.500 32.250 30.500 ;
        RECT 31.250 14.500 38.250 15.500 ;
        RECT 36.750 14.000 38.750 16.000 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 15.750 29.000 17.750 31.000 ;
        RECT 13.250 29.500 17.250 30.500 ;
        RECT 33.750 20.000 35.750 22.000 ;
        RECT 34.250 20.500 59.250 21.500 ;
        RECT 57.750 20.000 59.750 22.000 ;
        RECT 48.750 20.000 50.750 22.000 ;
        RECT 13.250 6.500 14.250 30.500 ;
        RECT 48.750 6.000 50.750 8.000 ;
        RECT 48.750 29.000 50.750 31.000 ;
        RECT 48.750 2.000 50.750 4.000 ;
        RECT 49.250 2.500 50.250 7.500 ;
        RECT 39.750 10.000 41.750 12.000 ;
        RECT 40.250 10.500 41.250 18.500 ;
        RECT 39.750 17.000 41.750 19.000 ;
        RECT 40.250 29.500 50.250 30.500 ;
        RECT 40.250 24.500 41.250 30.500 ;
        RECT 39.750 24.000 41.750 26.000 ;
        RECT 72.750 6.000 74.750 8.000 ;
        RECT 72.750 29.000 74.750 31.000 ;
        RECT 63.750 10.000 65.750 12.000 ;
        RECT 64.250 10.500 83.250 11.500 ;
        RECT 82.250 2.500 83.250 11.500 ;
        RECT 81.750 2.000 83.750 4.000 ;
        RECT 73.250 6.500 74.250 11.500 ;
        RECT 64.250 29.500 74.250 30.500 ;
        RECT 64.250 24.500 65.250 30.500 ;
        RECT 63.750 24.000 65.750 26.000 ;
  END
END DFQD1_2
MACRO DFQD1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFQD1_3 0 0 ; 
  SIZE 88.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN cp 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 10.500 11.250 15.500 ;
    END 
  END cp 
  PIN d 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 27.750 14.000 29.750 16.000 ;
        RECT 28.250 14.500 29.250 25.500 ;
        RECT 27.750 24.000 29.750 26.000 ;
    END 
  END d 
  PIN q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 78.750 6.000 80.750 8.000 ;
        RECT 78.750 29.000 80.750 31.000 ;
        RECT 79.250 6.500 80.250 30.500 ;
    END 
  END q 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 84.750 29.000 86.750 31.000 ;
        RECT 85.250 29.500 86.250 39.500 ;
        RECT 66.750 32.000 68.750 34.000 ;
        RECT 67.250 32.500 68.250 39.500 ;
        RECT 42.750 32.000 44.750 34.000 ;
        RECT 43.250 32.500 44.250 39.500 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 29.500 20.250 39.500 ;
        RECT 0.000 39.000 88.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 88.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 43.250 0.500 44.250 7.500 ;
        RECT 66.750 6.000 68.750 8.000 ;
        RECT 67.250 0.500 68.250 7.500 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 84.750 6.000 86.750 8.000 ;
        RECT 85.250 0.500 86.250 7.500 ;
        RECT 0.000 -1.000 88.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 88.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 12.750 2.000 14.750 4.000 ;
        RECT 13.250 2.500 14.250 7.500 ;
        RECT 15.750 29.000 17.750 31.000 ;
        RECT 13.250 29.500 17.250 30.500 ;
        RECT 54.750 6.000 56.750 8.000 ;
        RECT 54.750 29.000 56.750 31.000 ;
        RECT 55.250 2.500 56.250 7.500 ;
        RECT 54.750 2.000 56.750 4.000 ;
        RECT 69.750 20.000 71.750 22.000 ;
        RECT 70.250 20.500 71.250 25.500 ;
        RECT 55.250 24.500 71.250 25.500 ;
        RECT 55.250 24.500 56.250 30.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 2.500 32.250 7.500 ;
        RECT 30.750 2.000 32.750 4.000 ;
        RECT 31.250 6.500 32.250 30.500 ;
        RECT 31.250 24.500 47.250 25.500 ;
        RECT 45.750 24.000 47.750 26.000 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 33.750 17.000 35.750 19.000 ;
        RECT 34.250 17.500 59.250 18.500 ;
        RECT 57.750 17.000 59.750 19.000 ;
        RECT 51.750 14.000 53.750 16.000 ;
        RECT 52.250 14.500 53.250 18.500 ;
        RECT 1.250 6.500 2.250 18.500 ;
        RECT 1.250 17.500 23.250 18.500 ;
        RECT 21.750 17.000 23.750 19.000 ;
        RECT 48.750 6.000 50.750 8.000 ;
        RECT 48.750 29.000 50.750 31.000 ;
        RECT 48.750 20.000 50.750 22.000 ;
        RECT 49.250 20.500 50.250 30.500 ;
        RECT 49.250 6.500 50.250 15.500 ;
        RECT 43.250 14.500 50.250 15.500 ;
        RECT 42.750 14.000 44.750 16.000 ;
        RECT 72.750 6.000 74.750 8.000 ;
        RECT 72.750 29.000 74.750 31.000 ;
        RECT 63.750 10.000 65.750 12.000 ;
        RECT 64.250 10.500 77.250 11.500 ;
        RECT 75.750 10.000 77.750 12.000 ;
        RECT 73.250 10.500 74.250 30.500 ;
        RECT 73.250 6.500 74.250 21.500 ;
        RECT 72.750 20.000 74.750 22.000 ;
  END
END DFQD1_3
#--------EOF---------

MACRO FILL1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL1 0 0 ; 
  SIZE 2.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.000 39.000 2.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 2.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.000 -1.000 2.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 2.000 1.000 ;
    END 
  END vss 
END FILL1
#--------EOF---------

MACRO FILL2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL2 0 0 ; 
  SIZE 4.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.000 39.000 4.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 4.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.000 -1.000 4.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 4.000 1.000 ;
    END 
  END vss 
END FILL2
#--------EOF---------

MACRO FILL4
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL4 0 0 ; 
  SIZE 8.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.000 39.000 8.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 8.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.000 -1.000 8.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 8.000 1.000 ;
    END 
  END vss 
END FILL4
#--------EOF---------

MACRO FILL8
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILL8 0 0 ; 
  SIZE 16.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.000 39.000 16.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 16.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.000 -1.000 16.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 16.000 1.000 ;
    END 
  END vss 
END FILL8
#--------EOF---------

MACRO INVD1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVD1 0 0 ; 
  SIZE 10.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN i 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END i 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 6.500 2.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 0.000 39.000 10.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 10.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 0.000 -1.000 10.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 10.000 1.000 ;
    END 
  END vss 
END INVD1
#--------EOF---------

MACRO MUX2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1 0 0 ; 
  SIZE 46.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN i0 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 10.500 17.250 15.500 ;
    END 
  END i0 
  PIN i1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 10.500 11.250 15.500 ;
    END 
  END i1 
  PIN s 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 2.000 5.750 4.000 ;
        RECT 4.250 2.500 5.250 7.500 ;
    END 
  END s 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 43.250 6.500 44.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 37.250 29.500 38.250 39.500 ;
        RECT 0.000 39.000 46.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 46.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 36.750 6.000 38.750 8.000 ;
        RECT 37.250 0.500 38.250 7.500 ;
        RECT 0.000 -1.000 46.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 46.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 6.500 8.250 15.500 ;
        RECT 6.750 14.000 8.750 16.000 ;
        RECT 6.750 20.000 8.750 22.000 ;
        RECT 7.250 20.500 8.250 30.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 1.250 6.500 2.250 30.500 ;
        RECT 25.250 6.500 26.250 30.500 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 23.250 7.500 ;
        RECT 22.250 6.500 23.250 30.500 ;
        RECT 19.250 29.500 23.250 30.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 18.750 17.000 20.750 19.000 ;
        RECT 4.250 17.500 20.250 18.500 ;
        RECT 3.750 17.000 5.750 19.000 ;
        RECT 27.750 17.000 29.750 19.000 ;
        RECT 28.250 17.500 29.250 30.500 ;
        RECT 28.250 29.500 32.250 30.500 ;
        RECT 31.250 6.500 32.250 18.500 ;
        RECT 28.250 17.500 32.250 18.500 ;
  END
END MUX2D1
MACRO MUX2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1_1 0 0 ; 
  SIZE 46.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN i0 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 22.250 14.500 23.250 18.500 ;
    END 
  END i0 
  PIN i1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END i1 
  PIN s 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 2.000 11.750 4.000 ;
        RECT 10.250 2.500 11.250 7.500 ;
    END 
  END s 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 36.750 6.000 38.750 8.000 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 37.250 6.500 38.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 43.250 29.500 44.250 39.500 ;
        RECT 0.000 39.000 46.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 46.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 43.250 0.500 44.250 7.500 ;
        RECT 0.000 -1.000 46.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 46.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 6.500 8.250 30.500 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 6.500 23.250 7.500 ;
        RECT 22.250 6.500 23.250 11.500 ;
        RECT 22.250 10.500 35.250 11.500 ;
        RECT 34.250 2.500 35.250 11.500 ;
        RECT 34.250 2.500 41.250 3.500 ;
        RECT 39.750 2.000 41.750 4.000 ;
        RECT 13.250 6.500 14.250 30.500 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 20.250 30.500 ;
  END
END MUX2D1_1
MACRO MUX2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1_2 0 0 ; 
  SIZE 46.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN i0 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END i0 
  PIN i1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END i1 
  PIN s 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 22.250 14.500 23.250 18.500 ;
    END 
  END s 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 43.250 6.500 44.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 37.250 29.500 38.250 39.500 ;
        RECT 0.000 39.000 46.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 46.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 36.750 6.000 38.750 8.000 ;
        RECT 37.250 0.500 38.250 7.500 ;
        RECT 0.000 -1.000 46.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 46.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 20.250 30.500 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 25.250 6.500 26.250 30.500 ;
        RECT 1.250 6.500 2.250 30.500 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 6.500 8.250 30.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 30.750 2.000 32.750 4.000 ;
        RECT 31.250 2.500 32.250 7.500 ;
        RECT 31.250 6.500 32.250 30.500 ;
        RECT 30.750 24.000 32.750 26.000 ;
  END
END MUX2D1_2
MACRO MUX2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MUX2D1_3 0 0 ; 
  SIZE 46.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN i0 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END i0 
  PIN i1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 22.250 14.500 23.250 18.500 ;
    END 
  END i1 
  PIN s 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 27.750 2.000 29.750 4.000 ;
        RECT 28.250 2.500 29.250 7.500 ;
    END 
  END s 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 36.750 6.000 38.750 8.000 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 37.250 6.500 38.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 43.250 29.500 44.250 39.500 ;
        RECT 0.000 39.000 46.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 46.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 43.250 0.500 44.250 7.500 ;
        RECT 0.000 -1.000 46.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 46.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 20.250 30.500 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 6.500 17.250 7.500 ;
        RECT 16.250 2.500 17.250 7.500 ;
        RECT 16.250 2.500 23.250 3.500 ;
        RECT 22.250 2.500 23.250 11.500 ;
        RECT 22.250 10.500 35.250 11.500 ;
        RECT 34.250 2.500 35.250 11.500 ;
        RECT 34.250 2.500 41.250 3.500 ;
        RECT 39.750 2.000 41.750 4.000 ;
        RECT 13.250 6.500 14.250 30.500 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 6.500 8.250 30.500 ;
  END
END MUX2D1_3
#--------EOF---------

MACRO ND2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1 0 0 ; 
  SIZE 16.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 13.250 6.500 14.250 25.500 ;
        RECT 7.250 24.500 14.250 25.500 ;
        RECT 7.250 24.500 8.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 0.000 39.000 16.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 16.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 0.000 -1.000 16.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 16.000 1.000 ;
    END 
  END vss 
END ND2D1
MACRO ND2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1_1 0 0 ; 
  SIZE 16.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a2 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 1.250 6.500 2.250 25.500 ;
        RECT 1.250 24.500 8.250 25.500 ;
        RECT 7.250 24.500 8.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 0.000 39.000 16.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 16.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.000 -1.000 16.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 16.000 1.000 ;
    END 
  END vss 
END ND2D1_1
MACRO ND2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1_2 0 0 ; 
  SIZE 16.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 6.500 14.250 25.500 ;
        RECT 1.250 24.500 14.250 25.500 ;
        RECT 1.250 24.500 2.250 30.500 ;
        RECT 13.250 24.500 14.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 0.000 39.000 16.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 16.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 0.000 -1.000 16.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 16.000 1.000 ;
    END 
  END vss 
END ND2D1_2
MACRO ND2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND2D1_3 0 0 ; 
  SIZE 16.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 10.500 5.250 15.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a2 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 6.500 2.250 18.500 ;
        RECT 1.250 17.500 8.250 18.500 ;
        RECT 7.250 17.500 8.250 25.500 ;
        RECT 7.250 24.500 14.250 25.500 ;
        RECT 13.250 24.500 14.250 30.500 ;
        RECT 1.250 17.500 2.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 0.000 39.000 16.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 16.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.000 -1.000 16.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 16.000 1.000 ;
    END 
  END vss 
END ND2D1_3
#--------EOF---------

MACRO ND3D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1 0 0 ; 
  SIZE 28.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN a3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 22.250 14.500 23.250 18.500 ;
    END 
  END a3 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 13.250 6.500 14.250 25.500 ;
        RECT 13.250 24.500 20.250 25.500 ;
        RECT 19.250 24.500 20.250 30.500 ;
        RECT 7.250 24.500 14.250 25.500 ;
        RECT 7.250 24.500 8.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 0.000 39.000 28.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 28.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 0.000 -1.000 28.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 28.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 1.250 2.500 2.250 7.500 ;
        RECT 1.250 2.500 20.250 3.500 ;
        RECT 19.250 2.500 20.250 7.500 ;
  END
END ND3D1
MACRO ND3D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1_1 0 0 ; 
  SIZE 22.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a2 
  PIN a3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a3 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 7.250 6.500 20.250 7.500 ;
        RECT 7.250 6.500 8.250 30.500 ;
        RECT 7.250 24.500 20.250 25.500 ;
        RECT 19.250 24.500 20.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 0.000 39.000 22.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 22.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 0.000 -1.000 22.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 22.000 1.000 ;
    END 
  END vss 
END ND3D1_1
MACRO ND3D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1_2 0 0 ; 
  SIZE 28.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 22.250 14.500 23.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN a3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a3 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 20.250 18.500 ;
        RECT 13.250 17.500 20.250 18.500 ;
        RECT 13.250 17.500 14.250 25.500 ;
        RECT 7.250 24.500 14.250 25.500 ;
        RECT 7.250 24.500 8.250 30.500 ;
        RECT 19.250 17.500 20.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 0.000 39.000 28.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 28.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.000 -1.000 28.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 28.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 22.250 6.500 26.250 7.500 ;
        RECT 22.250 2.500 23.250 7.500 ;
        RECT 16.250 2.500 23.250 3.500 ;
        RECT 15.750 2.000 17.750 4.000 ;
        RECT 0.750 2.000 2.750 4.000 ;
        RECT 1.250 2.500 2.250 7.500 ;
  END
END ND3D1_2
MACRO ND3D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND3D1_3 0 0 ; 
  SIZE 28.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN a3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 22.250 14.500 23.250 18.500 ;
    END 
  END a3 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 13.250 6.500 14.250 30.500 ;
        RECT 1.250 24.500 14.250 25.500 ;
        RECT 1.250 24.500 2.250 30.500 ;
        RECT 13.250 29.500 20.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 0.000 39.000 28.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 28.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 0.000 -1.000 28.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 28.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 1.250 2.500 2.250 7.500 ;
        RECT 1.250 2.500 20.250 3.500 ;
        RECT 19.250 2.500 20.250 7.500 ;
  END
END ND3D1_3
#--------EOF---------

MACRO ND4D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1 0 0 ; 
  SIZE 34.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a2 
  PIN a3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a3 
  PIN a4 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 27.750 14.000 29.750 16.000 ;
        RECT 28.250 14.500 29.250 18.500 ;
    END 
  END a4 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 19.250 6.500 20.250 25.500 ;
        RECT 19.250 24.500 26.250 25.500 ;
        RECT 25.250 24.500 26.250 30.500 ;
        RECT 7.250 24.500 20.250 25.500 ;
        RECT 7.250 24.500 8.250 30.500 ;
        RECT 19.250 24.500 20.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 29.500 32.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 0.000 39.000 34.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 34.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 31.250 0.500 32.250 7.500 ;
        RECT 0.000 -1.000 34.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 34.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 25.250 2.500 26.250 7.500 ;
        RECT 1.250 2.500 26.250 3.500 ;
        RECT 1.250 2.500 2.250 7.500 ;
  END
END ND4D1
MACRO ND4D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1_1 0 0 ; 
  SIZE 34.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 27.750 14.000 29.750 16.000 ;
        RECT 28.250 14.500 29.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN a3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a3 
  PIN a4 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END a4 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 25.250 6.500 26.250 30.500 ;
        RECT 19.250 29.500 26.250 30.500 ;
        RECT 7.250 24.500 26.250 25.500 ;
        RECT 7.250 24.500 8.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 29.500 32.250 39.500 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 0.000 39.000 34.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 34.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 0.000 -1.000 34.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 34.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 1.250 6.500 17.250 7.500 ;
        RECT 16.250 6.500 17.250 11.500 ;
        RECT 16.250 10.500 23.250 11.500 ;
        RECT 22.250 2.500 23.250 11.500 ;
        RECT 22.250 2.500 32.250 3.500 ;
        RECT 31.250 2.500 32.250 7.500 ;
  END
END ND4D1_1
MACRO ND4D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1_2 0 0 ; 
  SIZE 28.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 22.250 14.500 23.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END a2 
  PIN a3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a3 
  PIN a4 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a4 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 25.250 6.500 26.250 25.500 ;
        RECT 19.250 24.500 26.250 25.500 ;
        RECT 19.250 24.500 20.250 30.500 ;
        RECT 7.250 24.500 20.250 25.500 ;
        RECT 7.250 24.500 8.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 0.000 39.000 28.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 28.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 0.000 -1.000 28.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 28.000 1.000 ;
    END 
  END vss 
END ND4D1_2
MACRO ND4D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ND4D1_3 0 0 ; 
  SIZE 34.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 27.750 14.000 29.750 16.000 ;
        RECT 28.250 14.500 29.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 22.250 14.500 23.250 18.500 ;
    END 
  END a2 
  PIN a3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a3 
  PIN a4 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a4 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 31.250 6.500 32.250 25.500 ;
        RECT 25.250 24.500 32.250 25.500 ;
        RECT 25.250 24.500 26.250 30.500 ;
        RECT 7.250 24.500 26.250 25.500 ;
        RECT 7.250 24.500 8.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 29.500 32.250 39.500 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 29.500 20.250 39.500 ;
        RECT 0.000 39.000 34.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 34.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.000 -1.000 34.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 34.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 16.250 6.500 20.250 7.500 ;
        RECT 16.250 6.500 17.250 11.500 ;
        RECT 1.250 10.500 17.250 11.500 ;
        RECT 1.250 6.500 2.250 11.500 ;
  END
END ND4D1_3
#--------EOF---------

MACRO NR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1 0 0 ; 
  SIZE 16.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a2 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 7.250 6.500 8.250 25.500 ;
        RECT 1.250 24.500 8.250 25.500 ;
        RECT 1.250 24.500 2.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 0.000 39.000 16.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 16.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.000 -1.000 16.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 16.000 1.000 ;
    END 
  END vss 
END NR2D1
MACRO NR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1_1 0 0 ; 
  SIZE 16.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 7.250 6.500 8.250 25.500 ;
        RECT 7.250 24.500 14.250 25.500 ;
        RECT 13.250 24.500 14.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 0.000 39.000 16.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 16.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 0.000 -1.000 16.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 16.000 1.000 ;
    END 
  END vss 
END NR2D1_1
MACRO NR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1_2 0 0 ; 
  SIZE 16.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a2 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 6.500 2.250 30.500 ;
        RECT 13.250 6.500 14.250 11.500 ;
        RECT 1.250 10.500 14.250 11.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 0.000 39.000 16.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 16.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 0.000 -1.000 16.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 16.000 1.000 ;
    END 
  END vss 
END NR2D1_2
MACRO NR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR2D1_3 0 0 ; 
  SIZE 16.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 6.500 14.250 30.500 ;
        RECT 1.250 6.500 2.250 11.500 ;
        RECT 1.250 10.500 14.250 11.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 0.000 39.000 16.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 16.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 0.000 -1.000 16.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 16.000 1.000 ;
    END 
  END vss 
END NR2D1_3
#--------EOF---------

MACRO NR3D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1 0 0 ; 
  SIZE 58.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 2.000 5.750 4.000 ;
        RECT 4.250 2.500 5.250 21.500 ;
        RECT 3.750 20.000 5.750 22.000 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 10.000 23.750 12.000 ;
        RECT 22.250 10.500 23.250 21.500 ;
        RECT 16.250 20.500 23.250 21.500 ;
        RECT 15.750 20.000 17.750 22.000 ;
    END 
  END a2 
  PIN a3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a3 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 6.500 11.250 7.500 ;
        RECT 10.250 6.500 11.250 11.500 ;
        RECT 10.250 10.500 20.250 11.500 ;
        RECT 19.250 6.500 20.250 11.500 ;
        RECT 7.250 6.500 8.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 43.250 29.500 44.250 39.500 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 29.500 32.250 39.500 ;
        RECT 0.000 39.000 58.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 58.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.000 -1.000 58.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 58.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 48.750 29.000 50.750 31.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 46.250 29.500 50.250 30.500 ;
        RECT 46.250 24.500 47.250 30.500 ;
        RECT 10.250 24.500 47.250 25.500 ;
        RECT 10.250 24.500 11.250 33.500 ;
        RECT 1.250 32.500 11.250 33.500 ;
        RECT 1.250 29.500 2.250 33.500 ;
        RECT 54.750 29.000 56.750 31.000 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 52.250 29.500 56.250 30.500 ;
        RECT 52.250 29.500 53.250 33.500 ;
        RECT 46.250 32.500 53.250 33.500 ;
        RECT 46.250 32.500 47.250 37.500 ;
        RECT 45.750 36.000 47.750 38.000 ;
        RECT 39.750 36.000 41.750 38.000 ;
        RECT 40.250 29.500 41.250 37.500 ;
        RECT 37.250 29.500 41.250 30.500 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 29.500 26.250 30.500 ;
  END
END NR3D1
MACRO NR3D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1_1 0 0 ; 
  SIZE 64.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 2.000 23.750 4.000 ;
        RECT 22.250 2.500 23.250 21.500 ;
        RECT 21.750 20.000 23.750 22.000 ;
    END 
  END a2 
  PIN a3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a3 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 6.500 11.250 7.500 ;
        RECT 10.250 6.500 11.250 11.500 ;
        RECT 10.250 10.500 20.250 11.500 ;
        RECT 19.250 6.500 20.250 11.500 ;
        RECT 7.250 6.500 8.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 48.750 29.000 50.750 31.000 ;
        RECT 49.250 29.500 50.250 39.500 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 37.250 29.500 38.250 39.500 ;
        RECT 0.000 39.000 64.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 64.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 0.000 -1.000 64.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 64.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 54.750 29.000 56.750 31.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 52.250 29.500 56.250 30.500 ;
        RECT 52.250 24.500 53.250 30.500 ;
        RECT 13.250 24.500 53.250 25.500 ;
        RECT 13.250 24.500 14.250 30.500 ;
        RECT 60.750 29.000 62.750 31.000 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 58.250 29.500 62.250 30.500 ;
        RECT 58.250 29.500 59.250 33.500 ;
        RECT 52.250 32.500 59.250 33.500 ;
        RECT 52.250 32.500 53.250 37.500 ;
        RECT 51.750 36.000 53.750 38.000 ;
        RECT 45.750 36.000 47.750 38.000 ;
        RECT 46.250 29.500 47.250 37.500 ;
        RECT 43.250 29.500 47.250 30.500 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 32.250 30.500 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 16.250 29.500 20.250 30.500 ;
        RECT 16.250 29.500 17.250 33.500 ;
        RECT 1.250 32.500 17.250 33.500 ;
        RECT 1.250 29.500 2.250 33.500 ;
  END
END NR3D1_1
MACRO NR3D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1_2 0 0 ; 
  SIZE 58.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 20.000 11.750 22.000 ;
        RECT 10.250 17.500 11.250 21.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 2.000 17.750 4.000 ;
        RECT 16.250 2.500 17.250 21.500 ;
        RECT 15.750 20.000 17.750 22.000 ;
    END 
  END a2 
  PIN a3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a3 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 1.250 6.500 5.250 7.500 ;
        RECT 4.250 6.500 5.250 11.500 ;
        RECT 4.250 10.500 14.250 11.500 ;
        RECT 13.250 6.500 14.250 11.500 ;
        RECT 7.250 10.500 8.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 43.250 29.500 44.250 39.500 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 29.500 32.250 39.500 ;
        RECT 0.000 39.000 58.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 58.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 0.000 -1.000 58.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 58.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 48.750 29.000 50.750 31.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 46.250 29.500 50.250 30.500 ;
        RECT 46.250 24.500 47.250 30.500 ;
        RECT 10.250 24.500 47.250 25.500 ;
        RECT 10.250 24.500 11.250 33.500 ;
        RECT 1.250 32.500 11.250 33.500 ;
        RECT 1.250 29.500 2.250 33.500 ;
        RECT 54.750 29.000 56.750 31.000 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 52.250 29.500 56.250 30.500 ;
        RECT 52.250 29.500 53.250 33.500 ;
        RECT 46.250 32.500 53.250 33.500 ;
        RECT 46.250 32.500 47.250 37.500 ;
        RECT 45.750 36.000 47.750 38.000 ;
        RECT 39.750 36.000 41.750 38.000 ;
        RECT 40.250 29.500 41.250 37.500 ;
        RECT 37.250 29.500 41.250 30.500 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 29.500 26.250 30.500 ;
  END
END NR3D1_2
MACRO NR3D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR3D1_3 0 0 ; 
  SIZE 58.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 10.000 23.750 12.000 ;
        RECT 22.250 10.500 23.250 21.500 ;
        RECT 16.250 20.500 23.250 21.500 ;
        RECT 15.750 20.000 17.750 22.000 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 20.000 26.750 22.000 ;
        RECT 25.250 20.500 53.250 21.500 ;
        RECT 51.750 20.000 53.750 22.000 ;
    END 
  END a2 
  PIN a3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END a3 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 16.250 6.500 20.250 7.500 ;
        RECT 16.250 6.500 17.250 11.500 ;
        RECT 7.250 10.500 17.250 11.500 ;
        RECT 7.250 6.500 8.250 11.500 ;
        RECT 13.250 10.500 14.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 43.250 29.500 44.250 39.500 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 29.500 32.250 39.500 ;
        RECT 0.000 39.000 58.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 58.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 0.000 -1.000 58.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 58.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 48.750 29.000 50.750 31.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 46.250 29.500 50.250 30.500 ;
        RECT 46.250 24.500 47.250 30.500 ;
        RECT 19.250 24.500 47.250 25.500 ;
        RECT 19.250 24.500 20.250 30.500 ;
        RECT 54.750 29.000 56.750 31.000 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 52.250 29.500 56.250 30.500 ;
        RECT 52.250 29.500 53.250 33.500 ;
        RECT 46.250 32.500 53.250 33.500 ;
        RECT 46.250 32.500 47.250 37.500 ;
        RECT 45.750 36.000 47.750 38.000 ;
        RECT 39.750 36.000 41.750 38.000 ;
        RECT 40.250 29.500 41.250 37.500 ;
        RECT 37.250 29.500 41.250 30.500 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 22.250 29.500 26.250 30.500 ;
        RECT 22.250 29.500 23.250 33.500 ;
        RECT 1.250 32.500 23.250 33.500 ;
        RECT 1.250 29.500 2.250 33.500 ;
  END
END NR3D1_3
#--------EOF---------

MACRO NR4D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR4D1 0 0 ; 
  SIZE 82.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 2.000 5.750 4.000 ;
        RECT 4.250 2.500 5.250 21.500 ;
        RECT 3.750 20.000 5.750 22.000 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 20.000 26.750 22.000 ;
        RECT 25.250 20.500 41.250 21.500 ;
        RECT 39.750 20.000 41.750 22.000 ;
    END 
  END a2 
  PIN a3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 48.750 20.000 50.750 22.000 ;
        RECT 49.250 20.500 77.250 21.500 ;
        RECT 75.750 20.000 77.750 22.000 ;
    END 
  END a3 
  PIN a4 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 27.750 14.000 29.750 16.000 ;
        RECT 28.250 14.500 29.250 18.500 ;
    END 
  END a4 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 22.250 6.500 26.250 7.500 ;
        RECT 22.250 6.500 23.250 11.500 ;
        RECT 7.250 10.500 23.250 11.500 ;
        RECT 7.250 6.500 8.250 11.500 ;
        RECT 7.250 10.500 8.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 66.750 29.000 68.750 31.000 ;
        RECT 67.250 29.500 68.250 39.500 ;
        RECT 54.750 29.000 56.750 31.000 ;
        RECT 55.250 29.500 56.250 39.500 ;
        RECT 0.000 39.000 82.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 82.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 31.250 0.500 32.250 7.500 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.000 -1.000 82.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 82.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 72.750 29.000 74.750 31.000 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 70.250 29.500 74.250 30.500 ;
        RECT 70.250 24.500 71.250 30.500 ;
        RECT 43.250 24.500 71.250 25.500 ;
        RECT 43.250 24.500 44.250 30.500 ;
        RECT 78.750 29.000 80.750 31.000 ;
        RECT 48.750 29.000 50.750 31.000 ;
        RECT 76.250 29.500 80.250 30.500 ;
        RECT 76.250 29.500 77.250 33.500 ;
        RECT 70.250 32.500 77.250 33.500 ;
        RECT 70.250 32.500 71.250 37.500 ;
        RECT 69.750 36.000 71.750 38.000 ;
        RECT 51.750 36.000 53.750 38.000 ;
        RECT 52.250 29.500 53.250 37.500 ;
        RECT 49.250 29.500 53.250 30.500 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 10.250 29.500 20.250 30.500 ;
        RECT 10.250 29.500 11.250 33.500 ;
        RECT 1.250 32.500 11.250 33.500 ;
        RECT 1.250 29.500 2.250 33.500 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 22.250 29.500 38.250 30.500 ;
        RECT 22.250 24.500 23.250 30.500 ;
        RECT 13.250 24.500 23.250 25.500 ;
        RECT 13.250 24.500 14.250 30.500 ;
  END
END NR4D1
MACRO NR4D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR4D1_1 0 0 ; 
  SIZE 76.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 20.000 20.750 22.000 ;
        RECT 19.250 20.500 35.250 21.500 ;
        RECT 33.750 20.000 35.750 22.000 ;
    END 
  END a2 
  PIN a3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 42.750 20.000 44.750 22.000 ;
        RECT 43.250 20.500 71.250 21.500 ;
        RECT 69.750 20.000 71.750 22.000 ;
    END 
  END a3 
  PIN a4 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 22.250 14.500 23.250 18.500 ;
    END 
  END a4 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 16.250 6.500 20.250 7.500 ;
        RECT 16.250 6.500 17.250 11.500 ;
        RECT 7.250 10.500 17.250 11.500 ;
        RECT 7.250 6.500 8.250 11.500 ;
        RECT 7.250 10.500 8.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 60.750 29.000 62.750 31.000 ;
        RECT 61.250 29.500 62.250 39.500 ;
        RECT 48.750 29.000 50.750 31.000 ;
        RECT 49.250 29.500 50.250 39.500 ;
        RECT 0.000 39.000 76.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 76.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 0.000 -1.000 76.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 76.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 66.750 29.000 68.750 31.000 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 64.250 29.500 68.250 30.500 ;
        RECT 64.250 24.500 65.250 30.500 ;
        RECT 37.250 24.500 65.250 25.500 ;
        RECT 37.250 24.500 38.250 30.500 ;
        RECT 72.750 29.000 74.750 31.000 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 70.250 29.500 74.250 30.500 ;
        RECT 70.250 29.500 71.250 33.500 ;
        RECT 64.250 32.500 71.250 33.500 ;
        RECT 64.250 32.500 65.250 37.500 ;
        RECT 63.750 36.000 65.750 38.000 ;
        RECT 45.750 36.000 47.750 38.000 ;
        RECT 46.250 29.500 47.250 37.500 ;
        RECT 43.250 29.500 47.250 30.500 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 10.250 29.500 32.250 30.500 ;
        RECT 10.250 29.500 11.250 33.500 ;
        RECT 1.250 32.500 11.250 33.500 ;
        RECT 1.250 29.500 2.250 33.500 ;
  END
END NR4D1_1
MACRO NR4D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NR4D1_2 0 0 ; 
  SIZE 82.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 27.750 2.000 29.750 4.000 ;
        RECT 28.250 2.500 29.250 37.500 ;
        RECT 22.250 36.500 29.250 37.500 ;
        RECT 21.750 36.000 23.750 38.000 ;
        RECT 27.750 36.000 29.750 38.000 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 2.000 5.750 4.000 ;
        RECT 4.250 2.500 5.250 21.500 ;
        RECT 3.750 20.000 5.750 22.000 ;
        RECT 4.250 20.500 23.250 21.500 ;
        RECT 21.750 20.000 23.750 22.000 ;
    END 
  END a2 
  PIN a3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 48.750 20.000 50.750 22.000 ;
        RECT 49.250 20.500 77.250 21.500 ;
        RECT 75.750 20.000 77.750 22.000 ;
    END 
  END a3 
  PIN a4 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a4 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 7.250 6.500 11.250 7.500 ;
        RECT 10.250 6.500 11.250 11.500 ;
        RECT 10.250 10.500 26.250 11.500 ;
        RECT 25.250 6.500 26.250 11.500 ;
        RECT 25.250 10.500 26.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 66.750 29.000 68.750 31.000 ;
        RECT 67.250 29.500 68.250 39.500 ;
        RECT 54.750 29.000 56.750 31.000 ;
        RECT 55.250 29.500 56.250 39.500 ;
        RECT 0.000 39.000 82.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 82.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 31.250 0.500 32.250 7.500 ;
        RECT 0.000 -1.000 82.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 82.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 72.750 29.000 74.750 31.000 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 70.250 29.500 74.250 30.500 ;
        RECT 70.250 24.500 71.250 30.500 ;
        RECT 43.250 24.500 71.250 25.500 ;
        RECT 43.250 24.500 44.250 30.500 ;
        RECT 78.750 29.000 80.750 31.000 ;
        RECT 48.750 29.000 50.750 31.000 ;
        RECT 76.250 29.500 80.250 30.500 ;
        RECT 76.250 29.500 77.250 33.500 ;
        RECT 70.250 32.500 77.250 33.500 ;
        RECT 70.250 32.500 71.250 37.500 ;
        RECT 69.750 36.000 71.750 38.000 ;
        RECT 51.750 36.000 53.750 38.000 ;
        RECT 52.250 29.500 53.250 37.500 ;
        RECT 49.250 29.500 53.250 30.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 1.250 29.500 20.250 30.500 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 29.500 38.250 30.500 ;
  END
END NR4D1_2
#--------EOF---------

MACRO OA21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1 0 0 ; 
  SIZE 34.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 27.750 14.000 29.750 16.000 ;
        RECT 28.250 14.500 29.250 18.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 17.000 11.750 19.000 ;
        RECT 10.250 17.500 11.250 21.500 ;
    END 
  END b 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 20.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 29.500 32.250 39.500 ;
        RECT 0.000 39.000 34.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 34.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.000 -1.000 34.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 34.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 22.250 6.500 26.250 7.500 ;
        RECT 22.250 2.500 23.250 7.500 ;
        RECT 16.250 2.500 23.250 3.500 ;
        RECT 15.750 2.000 17.750 4.000 ;
        RECT 0.750 2.000 2.750 4.000 ;
        RECT 1.250 2.500 2.250 7.500 ;
        RECT 6.750 2.000 8.750 4.000 ;
        RECT 7.250 2.500 8.250 30.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 31.250 6.500 32.250 21.500 ;
        RECT 22.250 20.500 32.250 21.500 ;
        RECT 22.250 20.500 23.250 33.500 ;
        RECT 16.250 32.500 23.250 33.500 ;
        RECT 16.250 14.500 17.250 33.500 ;
        RECT 10.250 14.500 17.250 15.500 ;
        RECT 10.250 6.500 11.250 15.500 ;
        RECT 7.250 6.500 11.250 7.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 1.250 29.500 5.250 30.500 ;
        RECT 4.250 29.500 5.250 33.500 ;
        RECT 4.250 32.500 11.250 33.500 ;
        RECT 10.250 32.500 11.250 37.500 ;
        RECT 9.750 36.000 11.750 38.000 ;
        RECT 24.750 36.000 26.750 38.000 ;
        RECT 25.250 29.500 26.250 37.500 ;
  END
END OA21D1
MACRO OA21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1_1 0 0 ; 
  SIZE 34.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END b 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 6.500 26.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 29.500 32.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 29.500 20.250 39.500 ;
        RECT 0.000 39.000 34.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 34.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 31.250 0.500 32.250 7.500 ;
        RECT 0.000 -1.000 34.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 34.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 13.250 6.500 14.250 25.500 ;
        RECT 7.250 24.500 14.250 25.500 ;
        RECT 7.250 24.500 8.250 30.500 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 19.250 2.500 20.250 7.500 ;
        RECT 7.250 2.500 20.250 3.500 ;
        RECT 7.250 2.500 8.250 7.500 ;
  END
END OA21D1_1
MACRO OA21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1_2 0 0 ; 
  SIZE 34.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 14.000 2.750 16.000 ;
        RECT 1.250 14.500 2.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 17.000 11.750 19.000 ;
        RECT 10.250 17.500 11.250 21.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 17.000 17.750 19.000 ;
        RECT 16.250 17.500 17.250 21.500 ;
    END 
  END b 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 6.500 29.250 7.500 ;
        RECT 28.250 6.500 29.250 30.500 ;
        RECT 25.250 29.500 29.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 29.500 32.250 39.500 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 0.000 39.000 34.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 34.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 31.250 0.500 32.250 7.500 ;
        RECT 0.000 -1.000 34.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 34.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 7.250 6.500 8.250 25.500 ;
        RECT 7.250 24.500 20.250 25.500 ;
        RECT 19.250 24.500 20.250 30.500 ;
        RECT 24.750 14.000 26.750 16.000 ;
        RECT 4.250 14.500 26.250 15.500 ;
        RECT 4.250 14.500 5.250 30.500 ;
        RECT 1.250 29.500 5.250 30.500 ;
        RECT 7.250 14.500 11.250 15.500 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 13.250 2.500 14.250 7.500 ;
        RECT 1.250 2.500 14.250 3.500 ;
        RECT 1.250 2.500 2.250 7.500 ;
  END
END OA21D1_2
MACRO OA21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21D1_3 0 0 ; 
  SIZE 34.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 17.000 17.750 19.000 ;
        RECT 16.250 17.500 17.250 21.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END b 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 6.500 26.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 29.500 32.250 39.500 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 0.000 39.000 34.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 34.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 31.250 0.500 32.250 7.500 ;
        RECT 0.000 -1.000 34.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 34.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 13.250 6.500 14.250 25.500 ;
        RECT 13.250 24.500 20.250 25.500 ;
        RECT 19.250 24.500 20.250 30.500 ;
        RECT 18.750 14.000 20.750 16.000 ;
        RECT 13.250 14.500 20.250 15.500 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 7.250 2.500 8.250 7.500 ;
        RECT 7.250 2.500 20.250 3.500 ;
        RECT 19.250 2.500 20.250 7.500 ;
  END
END OA21D1_3
#--------EOF---------

MACRO OAI21D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1 0 0 ; 
  SIZE 22.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END b 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 13.250 6.500 14.250 25.500 ;
        RECT 7.250 24.500 14.250 25.500 ;
        RECT 7.250 24.500 8.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 29.500 20.250 39.500 ;
        RECT 0.000 39.000 22.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 22.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 0.000 -1.000 22.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 22.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 7.250 2.500 8.250 7.500 ;
        RECT 7.250 2.500 20.250 3.500 ;
        RECT 19.250 2.500 20.250 7.500 ;
  END
END OAI21D1
MACRO OAI21D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1_1 0 0 ; 
  SIZE 22.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 16.250 14.500 17.250 18.500 ;
    END 
  END b 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 7.250 6.500 8.250 25.500 ;
        RECT 7.250 24.500 14.250 25.500 ;
        RECT 13.250 24.500 14.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 29.500 20.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 0.000 39.000 22.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 22.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 0.000 -1.000 22.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 22.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 13.250 2.500 14.250 7.500 ;
        RECT 1.250 2.500 14.250 3.500 ;
        RECT 1.250 2.500 2.250 7.500 ;
  END
END OAI21D1_1
MACRO OAI21D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1_2 0 0 ; 
  SIZE 28.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 22.250 14.500 23.250 18.500 ;
    END 
  END b 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 1.250 6.500 2.250 30.500 ;
        RECT 1.250 24.500 20.250 25.500 ;
        RECT 19.250 24.500 20.250 30.500 ;
        RECT 13.250 6.500 17.250 7.500 ;
        RECT 15.750 6.000 17.750 8.000 ;
        RECT 15.750 24.000 17.750 26.000 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 0.000 39.000 28.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 28.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 0.000 -1.000 28.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 28.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 7.250 2.500 8.250 7.500 ;
        RECT 7.250 2.500 20.250 3.500 ;
        RECT 19.250 2.500 20.250 7.500 ;
  END
END OAI21D1_2
MACRO OAI21D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21D1_3 0 0 ; 
  SIZE 28.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN b 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 22.250 14.500 23.250 18.500 ;
    END 
  END b 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 13.250 6.500 17.250 7.500 ;
        RECT 15.750 6.000 17.750 8.000 ;
        RECT 15.750 29.000 17.750 31.000 ;
        RECT 13.250 29.500 17.250 30.500 ;
        RECT 16.250 29.500 20.250 30.500 ;
        RECT 1.250 2.500 2.250 7.500 ;
        RECT 1.250 2.500 14.250 3.500 ;
        RECT 13.250 2.500 14.250 7.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 0.000 39.000 28.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 28.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 0.000 -1.000 28.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 28.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 7.250 6.500 8.250 11.500 ;
        RECT 7.250 10.500 20.250 11.500 ;
        RECT 19.250 6.500 20.250 11.500 ;
  END
END OAI21D1_3
#--------EOF---------

MACRO OR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1 0 0 ; 
  SIZE 22.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a2 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 20.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 0.000 39.000 22.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 22.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 0.000 -1.000 22.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 22.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 6.750 2.000 8.750 4.000 ;
        RECT 7.250 2.500 8.250 7.500 ;
        RECT 7.250 6.500 8.250 25.500 ;
        RECT 1.250 24.500 8.250 25.500 ;
        RECT 1.250 24.500 2.250 30.500 ;
  END
END OR2D1
MACRO OR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1_1 0 0 ; 
  SIZE 28.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 20.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 0.000 39.000 28.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 28.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 0.500 14.250 7.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 0.000 -1.000 28.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 28.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 7.250 6.500 8.250 25.500 ;
        RECT 7.250 24.500 14.250 25.500 ;
        RECT 13.250 24.500 14.250 30.500 ;
  END
END OR2D1_1
MACRO OR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1_2 0 0 ; 
  SIZE 28.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a2 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 20.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 29.500 14.250 39.500 ;
        RECT 0.000 39.000 28.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 28.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 0.000 -1.000 28.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 28.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 21.750 2.000 23.750 4.000 ;
        RECT 13.250 2.500 23.250 3.500 ;
        RECT 13.250 2.500 14.250 7.500 ;
        RECT 1.250 6.500 2.250 30.500 ;
  END
END OR2D1_2
MACRO OR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2D1_3 0 0 ; 
  SIZE 28.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 14.000 11.750 16.000 ;
        RECT 10.250 14.500 11.250 18.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 23.250 7.500 ;
        RECT 22.250 6.500 23.250 30.500 ;
        RECT 19.250 29.500 23.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 0.000 39.000 28.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 28.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 0.000 -1.000 28.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 28.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 15.750 29.000 17.750 31.000 ;
        RECT 13.250 29.500 17.250 30.500 ;
        RECT 13.250 6.500 14.250 30.500 ;
        RECT 1.250 6.500 2.250 11.500 ;
        RECT 1.250 10.500 14.250 11.500 ;
  END
END OR2D1_3
#--------EOF---------

MACRO TAPCELL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TAPCELL 0 0 ; 
  SIZE 14.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 2.500 28.500 4.500 30.500 ;
        RECT 3.000 29.000 4.000 39.500 ;
        RECT 5.500 28.500 7.500 30.500 ;
        RECT 6.000 29.000 7.000 39.500 ;
        RECT 8.500 28.500 10.500 30.500 ;
        RECT 9.000 29.000 10.000 39.500 ;
        RECT 0.000 39.000 14.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 14.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 2.500 6.500 4.500 8.500 ;
        RECT 3.000 0.500 4.000 8.000 ;
        RECT 5.500 6.500 7.500 8.500 ;
        RECT 6.000 0.500 7.000 8.000 ;
        RECT 8.500 6.500 10.500 8.500 ;
        RECT 9.000 0.500 10.000 8.000 ;
        RECT 0.000 -1.000 14.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 14.000 1.000 ;
    END 
  END vss 
END TAPCELL
#--------EOF---------

MACRO TIEH
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TIEH 0 0 ; 
  SIZE 10.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 1.250 29.500 5.250 30.500 ;
        RECT 4.250 29.500 5.250 33.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 0.000 39.000 10.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 10.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 0.000 -1.000 10.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 10.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 6.500 5.250 7.500 ;
        RECT 4.250 2.500 5.250 7.500 ;
        RECT 3.750 2.000 5.750 4.000 ;
  END
END TIEH
#--------EOF---------

MACRO TIEL
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TIEL 0 0 ; 
  SIZE 10.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 1.250 6.500 5.250 7.500 ;
        RECT 4.250 6.500 5.250 11.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 29.500 8.250 39.500 ;
        RECT 0.000 39.000 10.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 10.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 7.250 0.500 8.250 7.500 ;
        RECT 0.000 -1.000 10.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 10.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 3.750 20.000 5.750 22.000 ;
        RECT 4.250 20.500 5.250 30.500 ;
        RECT 1.250 29.500 5.250 30.500 ;
  END
END TIEL
#--------EOF---------

MACRO XNR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1 0 0 ; 
  SIZE 46.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 27.750 2.000 29.750 4.000 ;
        RECT 28.250 2.500 29.250 7.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 36.750 6.000 38.750 8.000 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 37.250 6.500 38.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 43.250 29.500 44.250 39.500 ;
        RECT 0.000 39.000 46.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 46.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 43.250 0.500 44.250 7.500 ;
        RECT 0.000 -1.000 46.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 46.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 6.500 23.250 7.500 ;
        RECT 22.250 6.500 23.250 15.500 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 7.250 6.500 8.250 30.500 ;
        RECT 22.250 14.500 23.250 37.500 ;
        RECT 21.750 36.000 23.750 38.000 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 20.250 30.500 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 30.750 2.000 32.750 4.000 ;
        RECT 31.250 2.500 32.250 18.500 ;
        RECT 25.250 17.500 32.250 18.500 ;
        RECT 24.750 17.000 26.750 19.000 ;
        RECT 12.750 17.000 14.750 19.000 ;
        RECT 13.250 6.500 14.250 18.500 ;
        RECT 13.250 17.500 14.250 30.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 6.500 35.250 7.500 ;
        RECT 34.250 6.500 35.250 21.500 ;
        RECT 25.250 20.500 35.250 21.500 ;
        RECT 24.750 20.000 26.750 22.000 ;
        RECT 15.750 20.000 17.750 22.000 ;
        RECT 16.250 14.500 17.250 21.500 ;
        RECT 15.750 14.000 17.750 16.000 ;
        RECT 31.250 20.500 32.250 30.500 ;
  END
END XNR2D1
MACRO XNR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1_1 0 0 ; 
  SIZE 46.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 27.750 24.000 29.750 26.000 ;
        RECT 10.250 24.500 29.250 25.500 ;
        RECT 9.750 24.000 11.750 26.000 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 17.000 23.750 19.000 ;
        RECT 22.250 17.500 26.250 18.500 ;
    END 
  END a2 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 36.750 6.000 38.750 8.000 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 37.250 6.500 38.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 43.250 29.500 44.250 39.500 ;
        RECT 0.000 39.000 46.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 46.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 43.250 0.500 44.250 7.500 ;
        RECT 0.000 -1.000 46.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 46.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 2.500 20.250 7.500 ;
        RECT 4.250 2.500 20.250 3.500 ;
        RECT 3.750 2.000 5.750 4.000 ;
        RECT 19.250 29.500 20.250 33.500 ;
        RECT 4.250 32.500 20.250 33.500 ;
        RECT 4.250 24.500 5.250 33.500 ;
        RECT 3.750 24.000 5.750 26.000 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 6.500 8.250 30.500 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 6.500 14.250 15.500 ;
        RECT 13.250 14.500 32.250 15.500 ;
        RECT 30.750 14.000 32.750 16.000 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 6.500 35.250 7.500 ;
        RECT 34.250 6.500 35.250 30.500 ;
        RECT 31.250 29.500 35.250 30.500 ;
        RECT 15.750 20.000 17.750 22.000 ;
        RECT 16.250 20.500 35.250 21.500 ;
  END
END XNR2D1_1
MACRO XNR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1_2 0 0 ; 
  SIZE 46.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 2.000 23.750 4.000 ;
        RECT 22.250 2.500 23.250 7.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 17.000 20.750 19.000 ;
        RECT 19.250 17.500 20.250 21.500 ;
    END 
  END a2 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 43.250 6.500 44.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 29.500 20.250 39.500 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 37.250 29.500 38.250 39.500 ;
        RECT 0.000 39.000 46.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 46.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 36.750 6.000 38.750 8.000 ;
        RECT 37.250 0.500 38.250 7.500 ;
        RECT 0.000 -1.000 46.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 46.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 6.500 17.250 7.500 ;
        RECT 16.250 6.500 17.250 11.500 ;
        RECT 16.250 10.500 29.250 11.500 ;
        RECT 27.750 10.000 29.750 12.000 ;
        RECT 13.250 6.500 14.250 30.500 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 31.250 6.500 32.250 15.500 ;
        RECT 16.250 14.500 32.250 15.500 ;
        RECT 16.250 14.500 17.250 33.500 ;
        RECT 10.250 32.500 17.250 33.500 ;
        RECT 10.250 14.500 11.250 33.500 ;
        RECT 4.250 14.500 11.250 15.500 ;
        RECT 4.250 6.500 5.250 15.500 ;
        RECT 1.250 6.500 5.250 7.500 ;
        RECT 31.250 14.500 32.250 30.500 ;
        RECT 1.250 29.500 11.250 30.500 ;
  END
END XNR2D1_2
MACRO XNR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNR2D1_3 0 0 ; 
  SIZE 46.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 2.000 23.750 4.000 ;
        RECT 22.250 2.500 26.250 3.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
    END 
  END a2 
  PIN zn 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 6.500 32.250 30.500 ;
    END 
  END zn 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 29.500 20.250 39.500 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 37.250 29.500 38.250 39.500 ;
        RECT 0.000 39.000 46.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 46.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 36.750 6.000 38.750 8.000 ;
        RECT 37.250 0.500 38.250 7.500 ;
        RECT 0.000 -1.000 46.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 46.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 6.500 17.250 7.500 ;
        RECT 16.250 6.500 17.250 11.500 ;
        RECT 16.250 10.500 29.250 11.500 ;
        RECT 28.250 2.500 29.250 11.500 ;
        RECT 28.250 2.500 35.250 3.500 ;
        RECT 33.750 2.000 35.750 4.000 ;
        RECT 13.250 6.500 14.250 30.500 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 34.250 6.500 35.250 37.500 ;
        RECT 33.750 36.000 35.750 38.000 ;
        RECT 3.750 36.000 5.750 38.000 ;
        RECT 4.250 6.500 5.250 37.500 ;
        RECT 1.250 6.500 5.250 7.500 ;
        RECT 40.250 29.500 44.250 30.500 ;
        RECT 1.250 29.500 5.250 30.500 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 16.250 6.500 17.250 33.500 ;
        RECT 10.250 32.500 17.250 33.500 ;
        RECT 10.250 6.500 11.250 33.500 ;
        RECT 7.250 6.500 11.250 7.500 ;
        RECT 7.250 29.500 11.250 30.500 ;
  END
END XNR2D1_3
#--------EOF---------

MACRO XOR2D1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1 0 0 ; 
  SIZE 46.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 9.750 17.000 11.750 19.000 ;
        RECT 10.250 17.500 11.250 25.500 ;
        RECT 10.250 24.500 29.250 25.500 ;
        RECT 27.750 24.000 29.750 26.000 ;
        RECT 15.750 24.000 17.750 26.000 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 22.250 10.500 23.250 15.500 ;
    END 
  END a2 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 36.750 6.000 38.750 8.000 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 37.250 6.500 38.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 43.250 29.500 44.250 39.500 ;
        RECT 0.000 39.000 46.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 46.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 43.250 0.500 44.250 7.500 ;
        RECT 0.000 -1.000 46.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 46.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 6.500 8.250 30.500 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 13.250 6.500 14.250 21.500 ;
        RECT 13.250 20.500 29.250 21.500 ;
        RECT 27.750 20.000 29.750 22.000 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 2.500 20.250 7.500 ;
        RECT 4.250 2.500 20.250 3.500 ;
        RECT 3.750 2.000 5.750 4.000 ;
        RECT 19.250 29.500 20.250 33.500 ;
        RECT 4.250 32.500 20.250 33.500 ;
        RECT 4.250 24.500 5.250 33.500 ;
        RECT 3.750 24.000 5.750 26.000 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 15.750 17.000 17.750 19.000 ;
        RECT 16.250 17.500 32.250 18.500 ;
        RECT 31.250 17.500 32.250 30.500 ;
        RECT 31.250 6.500 32.250 18.500 ;
  END
END XOR2D1
MACRO XOR2D1_1
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1_1 0 0 ; 
  SIZE 46.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 2.000 5.750 4.000 ;
        RECT 4.250 2.500 8.250 3.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 20.000 17.750 22.000 ;
        RECT 16.250 20.500 17.250 25.500 ;
    END 
  END a2 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 43.250 6.500 44.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 37.250 29.500 38.250 39.500 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 29.500 20.250 39.500 ;
        RECT 0.000 39.000 46.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 46.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 36.750 6.000 38.750 8.000 ;
        RECT 37.250 0.500 38.250 7.500 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 0.000 -1.000 46.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 46.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 1.250 6.500 17.250 7.500 ;
        RECT 16.250 6.500 17.250 11.500 ;
        RECT 16.250 10.500 32.250 11.500 ;
        RECT 31.250 6.500 32.250 11.500 ;
        RECT 1.250 6.500 2.250 30.500 ;
        RECT 31.250 10.500 32.250 30.500 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 6.500 8.250 11.500 ;
        RECT 7.250 10.500 14.250 11.500 ;
        RECT 13.250 10.500 14.250 15.500 ;
        RECT 13.250 14.500 29.250 15.500 ;
        RECT 27.750 14.000 29.750 16.000 ;
        RECT 7.250 10.500 8.250 30.500 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 12.750 17.000 14.750 19.000 ;
        RECT 13.250 17.500 26.250 18.500 ;
        RECT 24.750 17.000 26.750 19.000 ;
        RECT 27.750 6.000 29.750 8.000 ;
        RECT 25.250 6.500 29.250 7.500 ;
        RECT 9.750 17.000 11.750 19.000 ;
        RECT 10.250 17.500 11.250 37.500 ;
        RECT 4.250 36.500 11.250 37.500 ;
        RECT 3.750 36.000 5.750 38.000 ;
        RECT 25.250 17.500 26.250 30.500 ;
  END
END XOR2D1_1
MACRO XOR2D1_2
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1_2 0 0 ; 
  SIZE 46.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 2.000 5.750 4.000 ;
        RECT 4.250 2.500 8.250 3.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 15.750 20.000 17.750 22.000 ;
        RECT 16.250 20.500 17.250 25.500 ;
    END 
  END a2 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 30.750 6.000 32.750 8.000 ;
        RECT 30.750 29.000 32.750 31.000 ;
        RECT 31.250 6.500 32.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 37.250 29.500 38.250 39.500 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 29.500 20.250 39.500 ;
        RECT 0.000 39.000 46.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 46.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 36.750 6.000 38.750 8.000 ;
        RECT 37.250 0.500 38.250 7.500 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 19.250 0.500 20.250 7.500 ;
        RECT 0.000 -1.000 46.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 46.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 1.250 6.500 17.250 7.500 ;
        RECT 16.250 6.500 17.250 11.500 ;
        RECT 16.250 10.500 29.250 11.500 ;
        RECT 28.250 2.500 29.250 11.500 ;
        RECT 28.250 2.500 35.250 3.500 ;
        RECT 33.750 2.000 35.750 4.000 ;
        RECT 42.750 2.000 44.750 4.000 ;
        RECT 43.250 2.500 44.250 7.500 ;
        RECT 1.250 6.500 2.250 30.500 ;
        RECT 43.250 6.500 44.250 30.500 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 6.500 8.250 11.500 ;
        RECT 7.250 10.500 14.250 11.500 ;
        RECT 13.250 10.500 14.250 15.500 ;
        RECT 13.250 14.500 29.250 15.500 ;
        RECT 27.750 14.000 29.750 16.000 ;
        RECT 7.250 10.500 8.250 30.500 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 9.750 17.000 11.750 19.000 ;
        RECT 10.250 17.500 26.250 18.500 ;
        RECT 24.750 17.000 26.750 19.000 ;
        RECT 24.750 2.000 26.750 4.000 ;
        RECT 25.250 2.500 26.250 7.500 ;
        RECT 10.250 17.500 11.250 37.500 ;
        RECT 4.250 36.500 11.250 37.500 ;
        RECT 3.750 36.000 5.750 38.000 ;
        RECT 25.250 17.500 26.250 30.500 ;
  END
END XOR2D1_2
MACRO XOR2D1_3
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2D1_3 0 0 ; 
  SIZE 46.000 BY 40.000 ; 
  SYMMETRY X Y ; 
  SITE obscore ; 
  PIN a1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 27.750 2.000 29.750 4.000 ;
        RECT 28.250 2.500 29.250 7.500 ;
    END 
  END a1 
  PIN a2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 3.750 14.000 5.750 16.000 ;
        RECT 4.250 14.500 5.250 18.500 ;
    END 
  END a2 
  PIN z 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER ML1 ;
        RECT 36.750 6.000 38.750 8.000 ;
        RECT 36.750 29.000 38.750 31.000 ;
        RECT 37.250 6.500 38.250 30.500 ;
    END 
  END z 
  PIN vdd 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 29.000 26.750 31.000 ;
        RECT 25.250 29.500 26.250 39.500 ;
        RECT 0.750 29.000 2.750 31.000 ;
        RECT 1.250 29.500 2.250 39.500 ;
        RECT 42.750 29.000 44.750 31.000 ;
        RECT 43.250 29.500 44.250 39.500 ;
        RECT 0.000 39.000 46.000 41.000 ;
      LAYER ML2 ;
        RECT 0.000 39.000 46.000 41.000 ;
    END 
  END vdd 
  PIN vss 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER ML1 ;
        RECT 24.750 6.000 26.750 8.000 ;
        RECT 25.250 0.500 26.250 7.500 ;
        RECT 0.750 6.000 2.750 8.000 ;
        RECT 1.250 0.500 2.250 7.500 ;
        RECT 42.750 6.000 44.750 8.000 ;
        RECT 43.250 0.500 44.250 7.500 ;
        RECT 0.000 -1.000 46.000 1.000 ;
      LAYER ML2 ;
        RECT 0.000 -1.000 46.000 1.000 ;
    END 
  END vss 
  OBS
      LAYER ML1 ;
        RECT 18.750 6.000 20.750 8.000 ;
        RECT 18.750 29.000 20.750 31.000 ;
        RECT 19.250 6.500 20.250 30.500 ;
        RECT 12.750 6.000 14.750 8.000 ;
        RECT 12.750 29.000 14.750 31.000 ;
        RECT 13.250 6.500 17.250 7.500 ;
        RECT 16.250 2.500 17.250 7.500 ;
        RECT 16.250 2.500 23.250 3.500 ;
        RECT 22.250 2.500 23.250 11.500 ;
        RECT 22.250 10.500 35.250 11.500 ;
        RECT 34.250 2.500 35.250 11.500 ;
        RECT 34.250 2.500 41.250 3.500 ;
        RECT 39.750 2.000 41.750 4.000 ;
        RECT 13.250 6.500 14.250 30.500 ;
        RECT 6.750 6.000 8.750 8.000 ;
        RECT 6.750 29.000 8.750 31.000 ;
        RECT 7.250 6.500 8.250 30.500 ;
        RECT 7.250 29.500 11.250 30.500 ;
        RECT 10.250 29.500 11.250 33.500 ;
        RECT 10.250 32.500 23.250 33.500 ;
        RECT 22.250 14.500 23.250 33.500 ;
        RECT 21.750 14.000 23.750 16.000 ;
        RECT 7.250 24.500 8.250 30.500 ;
        RECT 22.250 32.500 23.250 37.500 ;
        RECT 21.750 36.000 23.750 38.000 ;
  END
END XOR2D1_3
#--------EOF---------


END LIBRARY
